module moduleName #(
    parameters NUM_NEURONS = 4
) (
    ports
);
    
endmodule